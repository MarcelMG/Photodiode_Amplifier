* ADA4350 Macro-model
* Function: Switched gain amplifier and ADC driver
*
* Revision History:
* Rev 2.1 May 2015-ZF
* Copyright 2015 by Analog Devices
* 
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spicemodels/license
* for License Statement. Use of this model indicates your acceptance
* of the terms and provisions in the License Staement.
*
* Tested on MultSIm, SiMetrix(NGSpice), PSpice
*
* Not modeled: Distortion, PSRR, Overload Recovery, Disable, CMRR
*             SPI interface
*
* Parameters modeled include:
*   Vos, Ibias, Input CM limits and Typ output voltge swing over full supply range,
*   Open Loop Gain & Phase, Slew Rate, Output current limits, Voltage & Current Noise over temp,
*   Capacitive load drive, Quiescent and dynamic supply currents,
*   Shut Down pin functionality where applicable,
*   Single supply & offset supply functionality.
*
* Model parameters represent +/- 5V supply specifications
*
* Parameter variations with supply are not modeled
*
* Node Assignments:
* Node names begin with the letter N and numeric nodes correspond to the ADA4350 pin numbers.
* Nodes designated with names correspond to ADA4350 pins with matching pin names
* Node P5 is not an actual ADA4350 pin. It is provided to enable all feedback path switching.
* Refeer to the ADA4350 datasheet for further information on this model
*
*
.Subckt ADA4350 N10 N11 VCC VEE VDD DGND N12 N13 P0 P1 P2 P3 P4 P5 N25 N26 N3 N2 N28 27 1 4 5 6 7 8 9
*
*
*
*** TIA, two amplifiers and three internal resistors ***
X1	N11	N10	VCC	VEE	N12	TIA
X2	N28	N2	VCC	VEE	N3	Amp
X3	30	29	VCC	VEE	N26	Amp
R1	N26	29	Rideal	500
R2	N3	29	Rideal	500
R3	30	N25	Rideal	500
I1	VDD	DGND	50e-6
*
*
*** 6 switch pairs ***
X4	VDD	P0	P0N	Trigger
S0	9	N12	P0	P0N	FBsw
S6	1	9	P0	P0N	Outsw
*
X5	VDD	P1	P1N	Trigger
S1	8	N12	P1	P1N	FBsw
S7	1	8	P1	P1N	Outsw
*
X6	VDD	P2	P2N	Trigger
S2	7	N12	P2	P2N	FBsw
S8	1	7	P2	P2N	Outsw
*
X7	VDD	P3	P3N	Trigger
S3	6	N13	P3	P3N	FBsw
S9	27	6	P3	P3N	Outsw
*
X8	VDD	P4	P4N	Trigger
S4	5	N13	P4	P4N	FBsw
S10	27	5	P4	P4N	Outsw
*
X9	VDD	P5	P5N	Trigger
S5	4	N13	P5	P5N	FBsw
S11	27	4	P5	P5N	Outsw
*
*
.model	Rideal	res(T_ABS=-273)
.model	FBsw	vswitch(Von=0.201,Voff=0.199,ron=150,roff=1e9)
.model	Outsw	vswitch(Von=0.201,Voff=0.199,ron=300,roff=1e9)
*
.ends Main
*
*
**********************************************
.Subckt Trigger VDD Trig TrigN
**********************************************
e1	2	1	VDD	0	0.2353
v1	1	0	0.42
e2	2	TrigN	4	0	1
R2	4	0	Rideal	1e3
C1	4	0	100e-12
V2	3	0	0.2
Sx	3	4	Trig	TrigN	DSwitch
*
.model	DSwitch	vswitch(Von=0.201,Voff=0.199,ron=0.001,roff=1e6)
.model	Rideal	res(T_ABS=-273)
*
.ends Trigger
*
*
*
**********************************************
.Subckt TIA 100 101 102 103 104
**********************************************
***Power Supplies***
Rz	102	1020	Rideal	1e-6
Ibias	1020	103	dc	0.5e-3
DzPS	98	1020	diode
Iquies	1020	98	dc	3.5e-3
S1	98	103	106	113	Switch
R1	102	99	Rideal	1e7
R2	99	103	Rideal	1e7
e1	111	110	102	110	1
e2	110	112	110	103	1
e3	110	0	99	0	1
*
*
***Inputs***
S2	1	100	106	113	Switch
S3	9	101	106	113	Switch
VOS	1	2	dc	15e-6
IbiasP	110	2	dc	0.25e-12
IbiasN	110	9	dc	0.25e-12
RinCMP	110	2	Rideal	100e6
RinCMN	9	110	Rideal	100e6
CinCMP	110	2	3e-12
CinCMN	9	110	3e-12
IOS	9	2	0.1e-12
RinDiff	9	2	Rideal	1000e3
CinDiff	9	2	2.5e-12
*
*
***Non-Inverting Input with Clamp***
g1	3	110	110	2	0.001
RInP	3	110	Rideal	1e3
RX1	40	3	Rideal	0.001
DInP	40	41	diode
DInN	42	40	diode
VinP	111	41	dc	1.66
VinN	42	112	dc	0.96
*
*
***Vnoise***
hVn	6	5	Vmeas1	707.10678
Vmeas1	20	110	DC	0
Vvn	21	110	dc	0.65
Dvn	21	20	DVnoisy
hVn1	6	7	Vmeas2	707.10678
Vmeas2	22	110	dc	0
Vvn1	23	110	dc	0.65
Dvn1	23	22	DVnoisy
*
*
***Inoise***
FnIN	9	110	Vmeas3	0.7071068
Vmeas3	51	110	dc	0
VnIN	50	110	dc	0.65
DnIN	50	51	DINnoisy
FnIN1	110	9	Vmeas4	0.7071068
Vmeas4	53	110	dc	0
VnIN1	52	110	dc	0.65
DnIN1	52	53	DINnoisy
*
FnIP	2	110	Vmeas5	0.7071068
Vmeas5	31	110	dc	0
VnIP	30	110	dc	0.65
DnIP	30	31	DIPnoisy
FnIP1	110	2	Vmeas6	0.7071068
Vmeas6	33	110	dc	0
VnIP1	32	110	dc	0.65
DnIP1	32	33	DIPnoisy
*
*
***CMRR***
RcmrrP	3	10	Rideal	1e12
RcmrrN	10	9	Rideal	1e12
g10	11	110	10	110	-1e-10
Lcmrr	11	12	1e-12
Rcmrr	12	110	Rideal	1e3
e4	5	3	11	110	1
*
*
***Power Down***
VPD	111	80	dc	2
VPD1	81	0	dc	1.5
RPD	111	106	Rideal	1e6
ePD	80	113	82	0	1
RDP1	82	0	Rideal	1e3
CPD	82	0	1e-10
S5	81	82	83	113	Switch
CDP1	83	0	1e-12
RPD2	106	83	1e6
*
*
***Feedback Pin***
*RF	105	104	Rideal	0.001
*
*
***VFB Stage***
g200	200	110	7	9	1
R200	200	110	Rideal	250
DzSlewP	201	200	DzSlewP
DzSlewN	201	110	DzSlewN
*
*
***1st Pole***
g210	210	110	200	110	4.8269e-6
R210	210	110	Rideal	1473.66e6
C210	210	110	1e-012
*
*
***Output Voltage Clamp-1***
RX2	60	210	Rideal	0.001
DzVoutP	61	60	DzVoutP
DzVoutN	60	62	DzVoutN
DVoutP	61	63	diode
DVoutN	64	62	diode
VoutP	65	63	dc	5.96
VoutN	64	66	dc	5.98
e60	65	110	111	110	1.0296
e61	66	110	112	110	1.0296
*
*
*** 11 frequency stages***
g220	220	110	210	110	0.001
R220	220	110	Rideal	1000
C220	220	110	0.234e-12
*
g230	230	110	220	110	0.001
R230	230	110	Rideal	1000
*
g240	240	110	230	110	0.001
R240	240	110	Rideal	1000
*
g245	245	110	240	110	0.001
R245	245	110	Rideal	1000
*
g250	250	110	245	110	0.001
R250	250	110	Rideal	1000
*
g255	255	110	250	110	0.001
R255	255	110	Rideal	1000
*
g260	260	110	255	110	0.001
R260	260	110	Rideal	1000
*
g265	265	110	260	110	0.001
R265	265	110	Rideal	1000
*
g270	270	110	265	110	0.001
R270	270	110	Rideal	1000
*
e280	280	110	270	110	1
R280	280	285	Rideal	10
L280	285	281	2.17e-9
C280	281	282	10.588e-12
R281	282	110	Rideal	10.048
*
e290	290	110	285	110	1
R290	290	292	Rideal	10
L290	290	291	0.362e-9
C290	291	292	17.51e-12
R291	292	110	Rideal	17.097
e295	295	110	292	110	1.585
*
*
***Output Stage***
g300	300	110	295	110	0.001
R300	300	110	Rideal	1000
e301	301	110	300	110	1
Rout	302	303	Rideal	 31
Lout	303	310	 13e-9
Cout	310	110	 10e-12
*
*
***Output Current Limit***
H1	301	304	Vsense1	100
Vsense1	301	302	dc	0
VIoutP	305	304	dc	3.836
VIoutN	304	306	dc	3.436
DIoutP	307	305	diode
DIoutN	306	307	diode
Rx3	307	300	Rideal	0.001
*
*
***Output Clamp-2***
VoutP1	111	73	dc	0.825
VoutN1	74	112	dc	0.785
DVoutP1	75	73	diode
DVoutN1	74	75	diode
RX4	75	310	Rideal	0.001
*
*
***Supply Currents***
FIoVcc	314	110	Vmeas8	1
Vmeas8	310	311	dc	0
R314	110	314	Rideal	1e9
DzOVcc	110	314	diode
DOVcc	102	314	diode
RX5	311	312	Rideal	0.001
FIoVee	315	110	Vmeas9	1
Vmeas9	312	313	dc	0
R315	315	110	Rideal	1e9
DzOVee	315	110	diode
DOVee	315	103	diode
*
*
***Output Switch***
S4	104	313	106	113	Switch
*
*
*** Common Models ***
.model	diode	d(bv=100)
.model	Switch	vswitch(Von=1.55,Voff=1.45,ron=0.001,roff=1e6)
.model	DzVoutP	D(BV=4.3)
.model	DzVoutN	D(BV=4.3)
.model	DzSlewP	D(BV=21.193)
.model	DzSlewN	D(BV=21.193)
.model	DVnoisy	D(IS=9.26e-16 KF=9.51e-16)
.model	DINnoisy	D(IS=3.81e-23 KF=0.00e0)
.model	DIPnoisy	D(IS=3.81e-23 KF=0.00e0)
.model	Rideal	res(T_ABS=-273)
*
.ends TIA
*
*
*
**********************************************
.Subckt Amp 100 101 102 103 104
**********************************************
***Power Supplies***
Rz	102	1020	Rideal	1e-6
Ibias	1020	103	dc	0.5e-3
DzPS	98	1020	diode
Iquies	1020	98	dc	3.5e-3
S1	98	103	106	113	Switch
R1	1020	99	Rideal	1e7
R2	99	103	Rideal	1e7
e1	111	110	1020	110	1
e2	110	112	110	103	1
e3	110	0	99	0	1
*
*
***Inputs***
S2	1	100	106	113	Switch
S3	9	101	106	113	Switch
VOS	1	2	dc	50e-6
IbiasP	110	2	dc	0.06e-6
IbiasN	110	9	dc	0.06e-6
RinCMP	110	2	Rideal	100e6
RinCMN	9	110	Rideal	100e6
CinCMP	110	2	2.4e-12
CinCMN	9	110	2.4e-12
IOS	9	2	0.06e-6
RinDiff	9	2	Rideal	100e3
CinDiff	9	2	0.6e-12
*
*
***Non-Inverting Input with Clamp***
g1	3	110	110	2	0.001
RInP	3	110	Rideal	1e3
RX1	40	3	Rideal	0.001
DInP	40	41	diode
DInN	42	40	diode
VinP	111	41	dc	1.66
VinN	42	112	dc	0.46
*
*
***Vnoise***
hVn	6	5	Vmeas1	707.10678
Vmeas1	20	110	DC	0
Vvn	21	110	dc	0.65
Dvn	21	20	DVnoisy
hVn1	6	7	Vmeas2	707.10678
Vmeas2	22	110	dc	0
Vvn1	23	110	dc	0.65
Dvn1	23	22	DVnoisy
*
*
***Inoise***
FnIN	9	110	Vmeas3	0.7071068
Vmeas3	51	110	dc	0
VnIN	50	110	dc	0.65
DnIN	50	51	DINnoisy
FnIN1	110	9	Vmeas4	0.7071068
Vmeas4	53	110	dc	0
VnIN1	52	110	dc	0.65
DnIN1	52	53	DINnoisy
*
FnIP	2	110	Vmeas5	0.7071068
Vmeas5	31	110	dc	0
VnIP	30	110	dc	0.65
DnIP	30	31	DIPnoisy
FnIP1	110	2	Vmeas6	0.7071068
Vmeas6	33	110	dc	0
VnIP1	32	110	dc	0.65
DnIP1	32	33	DIPnoisy
*
*
***CMRR***
RcmrrP	3	10	Rideal	1e12
RcmrrN	10	9	Rideal	1e12
g10	11	110	10	110	-1e-10
Lcmrr	11	12	1e-12
Rcmrr	12	110	Rideal	1e3
e4	5	3	11	110	1
*
*
***Power Down***
VPD	111	80	dc	0.8
VPD1	81	0	dc	0.1
RPD	111	106	Rideal	1e6
ePD	80	113	82	0	1
RDP1	82	0	Rideal	1e3
CPD	82	0	1e-10
S5	81	82	83	113	Switch
CDP1	83	0	1e-12
RPD2	106	83	1e6
*
*
***Feedback Pin***
*RF	105	104	Rideal	0.001
*
*
***VFB Stage***
g200	200	110	7	9	1
R200	200	110	Rideal	250
DzSlewP	201	200	DzSlewP
DzSlewN	201	110	DzSlewN
*
*
***1st Pole***
g210	210	110	200	110	2.2953e-6
R210	210	110	Rideal	1233.76e6
C210	210	110	1e-012
*
*
***Output Voltage Clamp-1***
RX2	60	210	Rideal	0.001
DzVoutP	61	60	DzVoutP
DzVoutN	60	62	DzVoutN
DVoutP	61	63	diode
DVoutN	64	62	diode
VoutP	65	63	dc	5.44
VoutN	64	66	dc	5.44
e60	65	110	111	110	1.098
e61	66	110	112	110	1.098
*
*
*** 11 frequency stages***
g220	220	110	210	110	0.001
R220	220	110	Rideal	1000
C220	220	110	1.179e-12
*
g230	230	110	220	110	0.001
R230	230	110	Rideal	1000
C230	230	110	0.042e-12
*
g240	240	110	230	110	0.001
R240	240	110	Rideal	1000
C240	240	110	0.029e-12
*
g245	245	110	240	110	0.001
R245	245	110	Rideal	1000
C245	245	110	0.029e-12
*
g250	250	110	245	110	0.001
R250	250	110	Rideal	1000
C250	250	110	0.029e-12
*
g255	255	110	250	110	0.001
R255	255	110	Rideal	1000
C255	255	110	0.029e-12
*
g260	260	110	255	110	0.001
R260	260	110	Rideal	1000
C260	260	110	0.029e-12
*
g265	265	110	260	110	0.001
R265	265	110	Rideal	1000
*
g270	270	110	265	110	0.001
R270	270	110	Rideal	1000
*
e280	280	110	270	110	1
R280	280	285	Rideal	10
L280	285	281	7.65e-9
C280	281	282	1635.136e-12
R281	282	110	Rideal	7.747
*
e290	290	110	285	110	1
R290	290	292	Rideal	10
L290	290	291	2.01e-9
C290	291	292	875.35e-12
R291	292	110	Rideal	26.289
e295	295	110	292	110	1.38
*
*
***Output Stage***
g300	300	110	295	110	0.001
R300	300	110	Rideal	1000
e301	301	110	300	110	1
Rout	302	303	Rideal	 49
Lout	303	310	 5e-9
Cout	310	110	 .4e-12
*
*
***Output Current Limit***
H1	301	304	Vsense1	100
Vsense1	301	302	dc	0
VIoutP	305	304	dc	6.936
VIoutN	304	306	dc	3.636
DIoutP	307	305	diode
DIoutN	306	307	diode
Rx3	307	300	Rideal	0.001
*
*
***Output Clamp-2***
VoutP1	111	73	dc	0.855
VoutN1	74	112	dc	0.855
DVoutP1	75	73	diode
DVoutN1	74	75	diode
RX4	75	310	Rideal	0.001
*
*
***Supply Currents***
FIoVcc	314	110	Vmeas8	1
Vmeas8	310	311	dc	0
R314	110	314	Rideal	1e9
DzOVcc	110	314	diode
DOVcc	102	314	diode
RX5	311	312	Rideal	0.001
FIoVee	315	110	Vmeas9	1
Vmeas9	312	313	dc	0
R315	315	110	Rideal	1e9
DzOVee	315	110	diode
DOVee	315	103	diode
*
*
***Output Switch***
S4	104	313	106	113	Switch
*
*
*** Common Models ***
.model	diode	d(bv=100)
.model	Switch	vswitch(Von=0.15,Voff=0.05,ron=0.001,roff=1e6)
.model	DzVoutP	D(BV=4.3)
.model	DzVoutN	D(BV=4.3)
.model	DzSlewP	D(BV=13.546)
.model	DzSlewN	D(BV=13.546)
.model	DVnoisy	D(IS=9.42e-16 KF=3.89e-16)
.model	DINnoisy	D(IS=4.62e-17 KF=0.00e0)
.model	DIPnoisy	D(IS=4.62e-17 KF=0.00e0)
.model	Rideal	res(T_ABS=-273)
*
.ends Amp
